library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instr_mem is
    port(
        --input
        addr_instr  : in std_logic_vector(31 downto 0);
        --output
        rd_instr    : out std_logic_vector(31 downto 0)
    );
end instr_mem;

architecture rtl of instr_mem is

    type romtype is array (64 downto 0) of std_logic_vector(31 downto 0);
    signal mem: romtype;

    begin

        --the program loads two matrix from the memory to the accelerator and saves the result from the accelerator

		mem(0) <= "0000000000000000000000010" & "0000011"; --lw x2, x0 + 0
		mem(1) <= "0000000100000000000000011" & "0000011"; --lw x3, x0 + 16
        mem(2) <= "000000010000" & "00010" & "001" & "00010" & "0011011"; --slli x2, x2, 16
		mem(3) <= "000000000000" & "00011" & "001" & "00011" & "0011011"; --slli x3, x3, 0
        mem(4) <= "0000000" & "00011" & "00010" & "110" & "00010" & "0110011"; --or x2, x2, x3

		mem(5) <= "0000001" & "00010" & "00000" & "000" & "00000" & "0100011"; --sw x2, x0 + 32
		mem(6) <= "000000100000" & "00000" & "00000000" & "1100000"; --ToAcc x0 + 32
		
        mem(7) <= "000000000100" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 4
        mem(8) <= "000000000101" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 5
        mem(9) <= "000000000110" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 6
        mem(10) <= "000000000111" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 7
        mem(11) <= "000000001000" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 8
        mem(12) <= "000000001001" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 9
        mem(13) <= "000000001010" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 10
        mem(14) <= "000000001011" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 11
        mem(15) <= "000000001100" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 12

        mem(16) <= "000000010100" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 20
        mem(17) <= "000000010101" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 21
        mem(18) <= "000000010110" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 22
        mem(19) <= "000000010111" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 23
        mem(20) <= "000000011000" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 24
        mem(21) <= "000000011001" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 25
        mem(22) <= "000000011010" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 26
        mem(23) <= "000000011011" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 27
        mem(24) <= "000000011100" & "00000" & "00000000" & "1100100"; --ToAccB x0 + 28

        mem(25) <= "0000001" & "00000" & "00000" & "000" & "00000" & "1101100"; --fromAccB x0 + 32
        mem(26) <= "0000001" & "00000" & "00000" & "000" & "00001" & "1101100"; --fromAccB x0 + 33
        mem(27) <= "0000001" & "00000" & "00000" & "000" & "00010" & "1101100"; --fromAccB x0 + 34
        mem(28) <= "0000001" & "00000" & "00000" & "000" & "00011" & "1101100"; --fromAccB x0 + 35
        mem(29) <= "0000001" & "00000" & "00000" & "000" & "00100" & "1101100"; --fromAccB x0 + 36
        mem(30) <= "0000001" & "00000" & "00000" & "000" & "00101" & "1101100"; --fromAccB x0 + 37
        mem(31) <= "0000001" & "00000" & "00000" & "000" & "00110" & "1101100"; --fromAccB x0 + 38
        mem(32) <= "0000001" & "00000" & "00000" & "000" & "00111" & "1101100"; --fromAccB x0 + 39
        mem(33) <= "0000001" & "00000" & "00000" & "000" & "01000" & "1101100"; --fromAccB x0 + 40

        mem(34) <= "0000001000000000000000011" & "0000011"; --lw x3, x0 + 32
        mem(35) <= "0000001001000000000000011" & "0000011"; --lw x3, x0 + 36
        mem(36) <= "0000001010000000000000011" & "0000011"; --lw x3, x0 + 40

        mem(37) <=  "0000000" & "00011" & "00010" & "110" & "00010" & "0110011"; --or x2, x2, x3
        mem(38) <= "00000000100000000000000000010011"; --addi x0, x0, 8
        mem(39) <= "00000000000000000000000000010011";
        mem(40) <= "00000000000000000000000000010011";
        mem(41) <= "00000000000000000000000000010011";
        mem(42) <= "00000000000000000000000000010011";
        mem(43) <= "00000000000000000000000000010011";
        mem(44) <= "00000000000000000000000000010011";
        mem(45) <= "00000000000000000000000000010011";
        mem(46) <= "00000000000000000000000000010011";
        mem(47) <= "00000000000000000000000000010011";
        mem(48) <= "00000000000000000000000000010011";
        mem(49) <= "00000000000000000000000000010011";
        mem(50) <= "00000000000000000000000000010011";
        mem(51) <= "00000000000000000000000000010011";
        mem(52) <= "00000000000000000000000000010011";
        mem(53) <= "00000000000000000000000000010011";
        mem(54) <= "00000000000000000000000000010011";
        mem(55) <= "00000000000000000000000000010011";
        mem(56) <= "00000000000000000000000000010011";
        mem(57) <= "00000000000000000000000000010011";
        mem(58) <= "00000000000000000000000000010011";
        mem(59) <= "00000000000000000000000000010011";
        mem(60) <= "00000000000000000000000000010011";
        mem(61) <= "00000000000000000000000000010011";
        mem(62) <= "00000000000000000000000000010011";
        mem(63) <= "00000000000000000000000000010011";
        mem(64) <= "00000000000000000000000000010011";      

        process(addr_instr,mem)begin
            rd_instr <= mem(to_integer(unsigned(addr_instr(31 downto 2))));
        end process;
    end rtl;
